# Translation by Martin Str�mberg <ams@ludd.luth.se>.
0.0:Install version %s, Copyright (C) 1998-2000 Jim Hall\n
0.1:Detta �r fri mjukvara, och du �r v�lkommen att redistribuera den\n
0.2:under s�rskilda vilkor; se filen COPYING f�r detaljer.\n
0.3:Install kommer med ABSOLUT INGEN GARANTI\n
0.4:Install-programmet avslutades framg�ngsrikt.
0.5:Det blev %u fel och %u icke-fatala varningar.\n
1.0:Tryck p� n�gon tangent f�r att forts�tta
1.1:Var �r installeringsfilerna? (att installera ifr�n?)
1.2:Var ska filerna installeras? (att installera till?)
2.0:nej
2.1:ja
2.2:Vill du installera detta disksetet? [jn]
2.3:Forts�tta installera denna disk? [jn]
2.4:Installera detta packetet? [jn]
3.0:Diskset: 
3.1:I top-niv�-install
3.2:Installerar serien: 
3.3:Packet: 
3.4:Kan inte hitta datafilerna f�r denna installdisk!
3.5:F�rdiginstallerat denna diskserie.
3.6:FEL!  Misslyckades att installera N�DV�NDIGT packet.
3.7:VARNING!  Misslyckades installera ICKE-N�DV�NDIGT packet.
3.8:Du har kanske fel installeringsfloppy i floppydriven.
3.9:Dubbelkolla att du har den r�tta disken och f�rs�k igen.
3.10:Om du ska installera andra diskserier, var v�nlig och stoppa in
3.11:disk #1 av n�sta serie i floppydriven nu.
4.0:ICKE-N�DV�NDIGT
4.1:N�DV�NDIGT
4.2:SKIPPAT
